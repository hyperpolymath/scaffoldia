// SPDX-License-Identifier: PMPL-1.0-or-later
//
// GitHub Pages Setup
// Enable and configure GitHub Pages in bulk

module github

import os
import json

// PagesSource represents where Pages should build from
pub enum PagesSource {
	root_main       // / on main branch
	docs_main       // /docs on main branch
	root_gh_pages   // / on gh-pages branch
	gh_pages_branch // gh-pages branch (legacy)
}

// PagesSetupParams contains parameters for Pages setup
pub struct PagesSetupParams {
pub:
	repo_owner string
	repo_name  string
	source     PagesSource
	cname      string  // Custom domain (optional)
	theme      string  // Jekyll theme (optional)
	dry_run    bool
}

// PagesSetupResult contains the result of Pages setup
pub struct PagesSetupResult {
pub:
	repo_path      string
	success        bool
	pages_enabled  bool
	pages_url      string
	message        string
}

// Convert PagesSource to API parameters
fn (source PagesSource) to_api_params() (string, string) {
	return match source {
		.root_main { 'main', '/' }
		.docs_main { 'main', '/docs' }
		.root_gh_pages { 'gh-pages', '/' }
		.gh_pages_branch { 'gh-pages', '/' }
	}
}

// Setup GitHub Pages for a repository
pub fn setup_pages(params PagesSetupParams) !PagesSetupResult {
	repo_full := '${params.repo_owner}/${params.repo_name}'

	if params.dry_run {
		return PagesSetupResult{
			repo_path: repo_full
			success: true
			pages_enabled: false
			pages_url: 'https://${params.repo_owner}.github.io/${params.repo_name}'
			message: '[DRY RUN] Would enable Pages'
		}
	}

	// Step 1: Check if Pages is already enabled
	println('  Checking Pages status...')
	check_result := os.execute('gh api "/repos/${repo_full}/pages" 2>/dev/null')

	if check_result.exit_code == 0 {
		// Pages already exists
		pages_url := os.execute('gh api "/repos/${repo_full}/pages" --jq .html_url 2>/dev/null').output.trim()
		return PagesSetupResult{
			repo_path: repo_full
			success: true
			pages_enabled: true
			pages_url: pages_url
			message: 'Pages already enabled at ${pages_url}'
		}
	}

	// Step 2: Enable Pages with specified source
	println('  Enabling Pages...')
	branch, path := params.source.to_api_params()

	// Create the pages site
	enable_cmd := 'gh api -X POST "/repos/${repo_full}/pages" -f source[branch]=${branch} -f source[path]=${path}'
	enable_result := os.execute(enable_cmd)

	if enable_result.exit_code != 0 {
		return PagesSetupResult{
			repo_path: repo_full
			success: false
			pages_enabled: false
			pages_url: ''
			message: 'Failed to enable Pages: ${enable_result.output}'
		}
	}

	// Step 3: Set custom domain if provided
	if params.cname != '' {
		println('  Setting custom domain...')
		cname_cmd := 'gh api -X PUT "/repos/${repo_full}/pages" -f cname=${params.cname}'
		os.execute(cname_cmd)
	}

	// Step 4: Get Pages URL
	pages_url := 'https://${params.repo_owner}.github.io/${params.repo_name}'

	return PagesSetupResult{
		repo_path: repo_full
		success: true
		pages_enabled: true
		pages_url: pages_url
		message: 'Pages enabled at ${pages_url}'
	}
}

// Check if Pages is enabled for a repository
pub fn check_pages_enabled(repo_owner string, repo_name string) bool {
	repo_full := '${repo_owner}/${repo_name}'
	result := os.execute('gh api "/repos/${repo_full}/pages" 2>/dev/null')
	return result.exit_code == 0
}

// Get Pages URL for a repository
pub fn get_pages_url(repo_owner string, repo_name string) string {
	repo_full := '${repo_owner}/${repo_name}'
	result := os.execute('gh api "/repos/${repo_full}/pages" --jq .html_url 2>/dev/null')
	if result.exit_code == 0 {
		return result.output.trim()
	}
	return ''
}

// Deploy default Jekyll site
pub fn deploy_jekyll_site(repo_path string, source PagesSource) !bool {
	// Determine target directory
	target_dir := match source {
		.docs_main {
			os.join_path(repo_path, 'docs')
		}
		else {
			repo_path
		}
	}

	// Create target directory
	os.mkdir_all(target_dir) or {
		return error('Failed to create target directory: ${err}')
	}

	// Create _config.yml
	config_path := os.join_path(target_dir, '_config.yml')
	config_content := 'theme: jekyll-theme-minimal
title: Repository Documentation
description: Automatically generated documentation site

# Build settings
markdown: kramdown
'

	os.write_file(config_path, config_content) or {
		return error('Failed to write _config.yml: ${err}')
	}

	// Create index.md
	index_path := os.join_path(target_dir, 'index.md')
	index_content := '# Documentation

Welcome to the documentation site!

## Contents

- [Getting Started](#getting-started)
- [API Reference](#api-reference)

## Getting Started

This site was automatically generated by repo-batcher.

## API Reference

See the [GitHub repository]({{ site.github.repository_url }}) for more information.
'

	os.write_file(index_path, index_content) or {
		return error('Failed to write index.md: ${err}')
	}

	return true
}

// Setup Pages for multiple repositories
pub fn setup_pages_batch(repos []string, source PagesSource, cname string, dry_run bool) []PagesSetupResult {
	mut results := []PagesSetupResult{}

	for repo in repos {
		// Parse owner/repo format
		parts := repo.split('/')
		if parts.len != 2 {
			results << PagesSetupResult{
				repo_path: repo
				success: false
				pages_enabled: false
				pages_url: ''
				message: 'Invalid repo format (expected owner/repo)'
			}
			continue
		}

		println('Setting up Pages for ${repo}...')
		result := setup_pages(PagesSetupParams{
			repo_owner: parts[0]
			repo_name: parts[1]
			source: source
			cname: cname
			theme: 'jekyll-theme-minimal'
			dry_run: dry_run
		}) or {
			PagesSetupResult{
				repo_path: repo
				success: false
				pages_enabled: false
				pages_url: ''
				message: 'Error: ${err}'
			}
		}
		results << result
		println('  ${result.message}')
	}

	return results
}

// Print Pages setup summary
pub fn print_pages_summary(results []PagesSetupResult) {
	mut success := 0
	mut already_enabled := 0
	mut failed := 0

	for result in results {
		if result.success {
			if result.message.contains('already enabled') {
				already_enabled++
			} else {
				success++
			}
		} else {
			failed++
		}
	}

	println('')
	println('=== Pages Setup Summary ===')
	println('Total repositories: ${results.len}')
	println('Successfully enabled: ${success}')
	println('Already enabled: ${already_enabled}')
	println('Failed: ${failed}')
	println('')

	// Show URLs for newly enabled pages
	if success > 0 {
		println('Newly enabled Pages sites:')
		for result in results {
			if result.success && !result.message.contains('already') {
				println('  ${result.repo_path} -> ${result.pages_url}')
			}
		}
		println('')
	}
}
